`timescale 1ns/100ps
module test_modADD(); 

logic clk;
logic [31:0] a,b,p,r;


ADDmod #(32)
ADDER(.A(a),.B(b),.P(p),.R(r));

always #0.5 clk = ~clk;

initial
begin
  clk='b0;
  
  a='b11111011100000000001111111110010;
  b='b11111011100000000001111100110010;
  p='b11111011100000000001111111110011;
  #1;
  a='b11111001111100001111000011110000;
  b='b11111001000000001111111100000000;
  p='b11111010000000000001111000011110;
  #1;
  a='b11110000111100001111000011110000;
  b='b11111011000000001111111100000000;
  p='b11111100000000000001111000011110;
  #1;
  a=32'b11100000111100001111000011110000;
  b=32'b1110111000000001111111100000000;
  p=32'b11110000000000000001111000011110;
  #1;
  a=32'b11000000111100001111000011110000;
  b=32'b11011111000000001111111100000000;
  p=32'b11100000000000000001111000011110;
  #3;
  $finish;
end

always@(posedge clk)
begin
  #0.5;
  if (r==32'b11111011100000000001111100110001)
    begin
    $display ("-------Testbench Result-------");
    $display ("----------pass first----------");
    end
  else
    $display ("---------failed first---------");
  
  #1;
  if (r==32'b11111000111100011101000111010010)
    $display ("----------pass second----------");
  else
    $display ("---------failed second---------");
  
  #1;
  if (r==32'b11101111111100011101000111010010)
    $display ("----------pass third----------");
  else
    $display ("---------failed third---------");
    
  #1;
  if (r==32'b1100111111100011101000111010010)
    $display ("----------pass fourth----------");
  else
    $display ("---------failed fourth---------");
    
  #1;
  if (r==32'b10111111111100011101000111010010)
    $display ("----------pass fifth----------");
  else
    $display ("---------failed fifth---------");
end
endmodule
